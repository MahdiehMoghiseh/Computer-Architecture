module ThirdROM(
  input [4:0] in3,
  output reg [5:0] out3
);
  always @(*) begin
    case (in3)
      5'b00001 : out3 = 6'b000000;
      5'b00010 : out3 = 6'b000001;
      5'b00011 : out3 = 6'b000010;
      5'b00100 : out3 = 6'b000110;
      5'b00101 : out3 = 6'b000111;
      5'b00110 : out3 = 6'b001100;

      5'b00111 : out3 = 6'b010000;
      5'b01000 : out3 = 6'b010001;
      5'b01001 : out3 = 6'b010010;
      5'b01010 : out3 = 6'b010110;
      5'b01011 : out3 = 6'b010111;
      5'b01100 : out3 = 6'b011100;

      5'b01101 : out3 = 6'b100000;
      5'b01110 : out3 = 6'b100001;
      5'b01111 : out3 = 6'b100010;
      5'b10000 : out3 = 6'b100110;
      5'b10001 : out3 = 6'b100111;
      5'b10010 : out3 = 6'b101100;

      5'b10011 : out3 = 6'b110000;
      5'b10100 : out3 = 6'b110001;
      5'b10101 : out3 = 6'b110010;
      5'b10110 : out3 = 6'b110110;
      5'b10111 : out3 = 6'b110111;
      5'b11000 : out3 = 6'b111100;
      default : out3 = 6'b010010;
    endcase
    
  end
endmodule

